`ifndef __APB_PKG_SV__
 `define __APB_PKG_SV__

package apb_pkg;
 `include "apb_drv.sv"
endpackage : apb_pkg

`endif // guard
